package toplevel_params is
  constant fu_LSU_dataw : integer := 32;
  constant fu_LSU_addrw : integer := 4;
  constant fu_INPUT_statusw : integer := 8;
  constant fu_OUTPUT_statusw : integer := 8;
end toplevel_params;
